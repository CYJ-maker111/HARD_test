module pills (
    input        clk,      // ʱ�����루1kHz��
    input        k0,       // pin 54 �� �ܿ��أ�1=������
    input        k1,       // ȫ������
    input        k2,       // ��ʼ����/��ͣ
    input        k4,       // pin 60 �� ��������ģʽ
    input        k5,       // pin 61 �� ѡ������ÿ��ƿ����������
    input        k6,       // pin 63 �� ѡ��������ƿ������
    input        k7,       // ����״̬����
    input        switch,   // �л�����

    output [6:0] LG1,      // ״̬��ʾ
    output reg [3:0] LG2,      // ��ǰƿҩƬ����λ
    output reg [3:0] LG3,      // ��ǰƿҩƬ��ʮλ
    output reg [3:0] LG4,      // ��װ��ƿ����λ
    output reg [3:0] LG5,      // ��װ��ƿ��ʮλ
    output reg [3:0] LG6,      // ��װ��ƿ����λ
    output       buzzer    // ������
);

// ========== �������� ==========
parameter S_IDLE    = 3'b000;  // ����״̬
parameter S_PAUSE   = 3'b001;  // ��ͣ״̬��Ĭ��״̬��
parameter S_SETUP   = 3'b010;  // ����״̬
parameter S_RUN     = 3'b011;  // ����״̬
parameter S_ERROR   = 3'b100;  // ����״̬

// �߶�����ܱ��루��������
parameter SEG_S = 7'b1101101;  // S
parameter SEG_C = 7'b0111001;  // C
parameter SEG_P = 7'b1110011;  // P
parameter SEG_E = 7'b1111001;  // E
parameter SEG_BLANK = 7'b1111111;

// ������ģʽ
parameter BEEP_COMPLETE = 2'b00;   // �����ʾ��
parameter BEEP_ALARM    = 2'b01;   // ������
parameter BEEP_ALARM_FAST = 2'b10; // ���پ�����������״̬��

// ========== �Ĵ������� ==========
reg [2:0] state;           // ��չ״̬λ��3λ
reg beep_enable;           // ������ʹ�ܿ���
reg finished;              // ��ɱ�־

// ���ؼ��
reg switch_last;          // switch���ؼ��

// ��ʾֵ
reg [6:0] seg_state;

// ������Ƶ�����ɣ�500Hz��
reg [1:0] tone_counter;   // 2λ��������������500Hz
reg beep_tone;
reg [1:0] beep_mode;      // ������ģʽ
reg alarm_enable;         // ������ʹ�ܿ��ƣ�����/�رվ������ࣩ

reg [9:0] lighting_counter;// Ƶ����ʱ��
reg light_state;
reg [7:0] alarm_counter;  // ��������ʱ��

// ���ò��� - ʹ��BCD��ֱ�Ӵ洢
reg [3:0] total_hundreds, total_tens, total_ones;    // ��ƿ��BCD��
reg [3:0] pills_tens, pills_ones;                    // ÿƿҩƬ��BCD��

// ����״̬�Ĵ��� - ʹ��BCD��ֱ�Ӵ洢
reg [3:0] current_pills_tens, current_pills_ones;    // ��ǰƿҩƬ��BCD��
reg [3:0] done_hundreds, done_tens, done_ones;       // ��װ��ƿ��BCD��
reg [9:0] timer;               // 1���ʱ��
reg [11:0] beep_timer;         // ��������ʱ����12λ�����4�룩

// ����ѡ���־
reg setting_pills;  // 1:��������ÿƿҩƬ��
reg setting_total;  // 1:����������ƿ��

// ����״̬��־
reg error_flag;     // ����״̬��־

// ========== ����߼� ==========
// ���ؼ��
wire switch_rise;
assign switch_rise = switch && !switch_last;

// ========== ��Ƶ�� ============

always @(posedge clk) begin

    if(lighting_counter == 10'd999) begin
        lighting_counter <= 1'b0;
        if(light_state == 1'b1)
            light_state <= 1'b0;
        else
            light_state <= 1'b1;
    end
    else
        lighting_counter <= lighting_counter + 1'b1;    

end

// ========== ��״̬�� ==========
always @(posedge clk) begin
    // ������һ��״̬���ڱ��ؼ��
    switch_last <= switch;
    
    // ��������ʱ������
    if (beep_mode == BEEP_ALARM || beep_mode == BEEP_ALARM_FAST) begin
        if (alarm_counter == 8'd0) begin
            alarm_enable <= ~alarm_enable;  // �л��������Ŀ���/�ر�״̬
            
            // ���ò�ͬ�������Ľ���
            if (beep_mode == BEEP_ALARM) begin
                // ��׼��������ÿ����1�Σ���500ms����500ms��
                if (alarm_enable == 1'b1) begin
                    alarm_counter <= 8'd250; // 500ms����
                end else begin
                    alarm_counter <= 8'd250; // 500ms�ر�
                end
            end else begin
                // ���پ�����������״̬����ÿ����2�Σ���250ms����250ms��
                if (alarm_enable == 1'b1) begin
                    alarm_counter <= 8'd125; // 250ms����
                end else begin
                    alarm_counter <= 8'd125; // 250ms�ر�
                end
            end
        end else begin
            alarm_counter <= alarm_counter - 8'd1;
        end
    end else begin
        alarm_enable <= 1'b0;
        alarm_counter <= 8'd0;
    end
    
    // �ܿ��ؿ���
    if (!k0) begin
        state <= S_IDLE;
        // �������мĴ���
        current_pills_tens <= 4'b0000;
        current_pills_ones <= 4'b0000;
        done_hundreds <= 4'b0000;
        done_tens <= 4'b0000;
        done_ones <= 4'b0000;
        timer <= 10'b0000000000;
        beep_timer <= 12'b000000000000;
        beep_enable <= 1'b0;
        finished <= 1'b0;
        setting_pills <= 1'b0;
        setting_total <= 1'b0;
        error_flag <= 1'b0;
        beep_mode <= BEEP_COMPLETE;
        alarm_enable <= 1'b0;
        alarm_counter <= 8'd0;
        
        // Ĭ�����ã���ƿ��2��ÿƿ10Ƭ
        total_hundreds <= 4'b0000;
        total_tens <= 4'b0000;
        total_ones <= 4'b0010;  // 2
        
        pills_tens <= 4'b0001;  // ʮλ1
        pills_ones <= 4'b0000;  // ��λ0
    end
    // ���㰴ť
    else if (k1) begin
        current_pills_tens <= 4'b0000;
        current_pills_ones <= 4'b0000;
        done_hundreds <= 4'b0000;
        done_tens <= 4'b0000;
        done_ones <= 4'b0000;
        timer <= 10'b0000000000;
        beep_timer <= 12'b000000000000;
        if (!error_flag) begin  // ������ڴ���״̬�������������
            beep_enable <= 1'b0;
            beep_mode <= BEEP_COMPLETE;
            alarm_enable <= 1'b0;
            alarm_counter <= 8'd0;
        end
        finished <= 1'b0;
        // ע�⣺����������־����Ҫ�ֶ��������״̬
    end
    else begin
        // ��������ʱ���ƣ����������ʾ����Ч��
        if (beep_enable && beep_mode == BEEP_COMPLETE) begin
            // ����Ƿ�ȫ��װ��
            // BCD�Ƚ��߼����ȱȽϰ�λ���ٱȽ�ʮλ�����Ƚϸ�λ
            if ((done_hundreds > total_hundreds) ||
                (done_hundreds == total_hundreds && done_tens > total_tens) ||
                (done_hundreds == total_hundreds && done_tens == total_tens && done_ones >= total_ones)) begin
                // ȫ��װ�꣺����4��
                if (beep_timer < 12'b111110100000) begin  // 4000
                    beep_timer <= beep_timer + 12'b000000000001;
                end else begin
                    beep_enable <= 1'b0;
                    beep_timer <= 12'b000000000000;
                    finished <= 1'b1;
                end
            end else begin
                // װ��һƿ������30ms
                if (beep_timer < 12'b000000011110) begin  // 30
                    beep_timer <= beep_timer + 12'b000000000001;
                end else begin
                    beep_enable <= 1'b0;
                    beep_timer <= 12'b000000000000;
                end
            end
        end
        
        case (state)
            S_IDLE: begin
                if (k0) begin
                    // ����Ĭ�Ͻ�����ͣ״̬
                    state <= S_PAUSE;
                    // ��������״̬
                    current_pills_tens <= 4'b0000;
                    current_pills_ones <= 4'b0000;
                    done_hundreds <= 4'b0000;
                    done_tens <= 4'b0000;
                    done_ones <= 4'b0000;
                    finished <= 1'b0;
                    setting_pills <= 1'b0;
                    setting_total <= 1'b0;
                    error_flag <= 1'b0;
                    beep_mode <= BEEP_COMPLETE;
                    alarm_enable <= 1'b0;
                    alarm_counter <= 8'd0;
                end
            end
            
            S_PAUSE: begin
                // ������״̬����
                if (k7) begin
                    state <= S_ERROR;
                    error_flag <= 1'b1;
                    beep_mode <= BEEP_ALARM_FAST;  // �������״̬�����ÿ��پ�����
                    beep_enable <= 1'b1;          // ���÷�����
                    alarm_enable <= 1'b1;         // ��ʼ����
                end
                // ��������ģʽ - ��k4Ϊ1ʱ
                else if (k4) begin
                    state <= S_SETUP;
                    setting_pills <= 1'b0;
                    setting_total <= 1'b0;
                end
                // ��ʼ���� - k2Ϊ1ʱ��������״̬
                else if (k2) begin
                    state <= S_RUN;
                end
            end
            
            S_SETUP: begin
                // ������״̬����
                if (k7) begin
                    state <= S_ERROR;
                    error_flag <= 1'b1;
                    beep_mode <= BEEP_ALARM_FAST;  // �������״̬�����ÿ��پ�����
                    beep_enable <= 1'b1;          // ���÷�����
                    alarm_enable <= 1'b1;         // ��ʼ����
                end
                // �˳�����ģʽ - ��k4Ϊ0ʱ�ص���ͣ״̬
                else if (!k4) begin
                    state <= S_PAUSE;
                end
                else begin
                    // ����ѡ��
                    if (k5) begin
                        setting_pills <= 1'b1;
                        setting_total <= 1'b0;
                    end
                    else if (k6) begin
                        setting_total <= 1'b1;
                        setting_pills <= 1'b0;
                    end
                    
                    // �л�����ֵ - switch�����ش���
                    if (switch_rise) begin
                        if (setting_pills) begin
                            // ����ÿƿҩƬ����10��20��50��10
                            if (pills_tens == 4'b0001 && pills_ones == 4'b0000) begin // 10
                                pills_tens <= 4'b0010; // 20
                                pills_ones <= 4'b0000;
                            end
                            else if (pills_tens == 4'b0010 && pills_ones == 4'b0000) begin // 20
                                pills_tens <= 4'b0101; // 50
                                pills_ones <= 4'b0000;
                            end
                            else begin // 50������
                                pills_tens <= 4'b0001; // 10
                                pills_ones <= 4'b0000;
                            end
                        end
                        else if (setting_total) begin
                            // ������ƿ����2��10��50��100��2
                            if (total_hundreds == 4'b0000 && total_tens == 4'b0000 && total_ones == 4'b0010) begin // 2
                                total_hundreds <= 4'b0000;
                                total_tens <= 4'b0001; // 10
                                total_ones <= 4'b0000;
                            end
                            else if (total_hundreds == 4'b0000 && total_tens == 4'b0001 && total_ones == 4'b0000) begin // 10
                                total_hundreds <= 4'b0000;
                                total_tens <= 4'b0101; // 50
                                total_ones <= 4'b0000;
                            end
                            else if (total_hundreds == 4'b0000 && total_tens == 4'b0101 && total_ones == 4'b0000) begin // 50
                                total_hundreds <= 4'b0001; // 100
                                total_tens <= 4'b0000;
                                total_ones <= 4'b0000;
                            end
                            else begin // 100������
                                total_hundreds <= 4'b0000;
                                total_tens <= 4'b0000;
                                total_ones <= 4'b0010; // 2
                            end
                        end
                    end
                end
            end
            
            S_RUN: begin
                // ������״̬����
                if (k7) begin
                    state <= S_ERROR;
                    error_flag <= 1'b1;
                    beep_mode <= BEEP_ALARM_FAST;  // �������״̬�����ÿ��پ�����
                    beep_enable <= 1'b1;          // ���÷�����
                    alarm_enable <= 1'b1;         // ��ʼ����
                end
                // ��ͣ���ص���ͣ״̬��- k2Ϊ0ʱ��ͣ
                else if (!k2) begin
                    state <= S_PAUSE;
                end
                // ����Ƿ�ȫ��װ����δ��ɷ���
                else if (((done_hundreds > total_hundreds) ||
                         (done_hundreds == total_hundreds && done_tens > total_tens) ||
                         (done_hundreds == total_hundreds && done_tens == total_tens && done_ones >= total_ones)) && !finished) begin
                    if (!beep_enable) begin
                        beep_enable <= 1'b1;
                        beep_mode <= BEEP_COMPLETE;  // ʹ�������ʾ��ģʽ
                        beep_timer <= 12'b000000000000;
                    end
                end
                // ����װƿ - ����Ƿ�δ�������ƿ��
                else if (!((done_hundreds > total_hundreds) ||
                          (done_hundreds == total_hundreds && done_tens > total_tens) ||
                          (done_hundreds == total_hundreds && done_tens == total_tens && done_ones >= total_ones))) begin
                    // 1��װһƬ
                    if (timer < 10'b1111100111) begin  // 999
                        timer <= timer + 10'b0000000001;
                    end
                    else begin
                        timer <= 10'b0000000000;  // 1�뵽
                        
                        // ��鵱ǰƿ�Ƿ�����
                        // �Ƚϵ�ǰҩƬ���Ƿ�С������ֵ
                        if ((current_pills_tens < pills_tens) || 
                            (current_pills_tens == pills_tens && current_pills_ones < pills_ones)) begin
                            // ��ǰƿδ����ҩƬ����1��BCD�ӷ���
                            if (current_pills_ones == 4'b1001) begin  // ��λΪ9
                                current_pills_ones <= 4'b0000;
                                current_pills_tens <= current_pills_tens + 4'b0001;
                            end else begin
                                current_pills_ones <= current_pills_ones + 4'b0001;
                            end
                        end
                        else begin
                            // ��ǰƿ����
                            current_pills_tens <= 4'b0000;
                            current_pills_ones <= 4'b0000;
                            
                            // ��װƿ����1��BCD�ӷ���
                            if (done_ones == 4'b1001) begin  // ��λΪ9
                                done_ones <= 4'b0000;
                                if (done_tens == 4'b1001) begin  // ʮλΪ9
                                    done_tens <= 4'b0000;
                                    done_hundreds <= done_hundreds + 4'b0001;
                                end else begin
                                    done_tens <= done_tens + 4'b0001;
                                end
                            end else begin
                                done_ones <= done_ones + 4'b0001;
                            end
                            
                            // ����һ����30ms��
                            beep_enable <= 1'b1;
                            beep_mode <= BEEP_COMPLETE;  // ʹ�������ʾ��ģʽ
                            beep_timer <= 12'b000000000000;
                        end
                    end
                end
            end
            
            S_ERROR: begin
                // ����״̬�����в�����ͣ
                // ֻ��k7Ϊ0ʱ�����˳�����״̬
                if (!k7) begin
                    error_flag <= 1'b0;   // ��������־
                    state <= S_PAUSE;     // �ص���ͣ״̬
                    beep_mode <= BEEP_COMPLETE; // �ָ�Ĭ�Ϸ���ģʽ
                    beep_enable <= 1'b0;  // �رշ�����
                    alarm_enable <= 1'b0; // �رվ�����
                    alarm_counter <= 8'd0; // ���ü�����
                end
                // ����״̬�³���������
            end
        endcase
    end
end

// ========== ���������߼� ==========
always @(posedge clk) begin
    if (tone_counter == 2'b01) begin
        tone_counter <= 2'b00;
        beep_tone <= ~beep_tone;  // ÿ2�����ڷ�תһ�� = 500Hz
    end else begin
        tone_counter <= tone_counter + 2'b01;
    end
end

// ========== ��ʾ�߼� ==========
always @(posedge clk) begin
    // ״̬��ʾ
    case (state)
        S_SETUP: seg_state <= SEG_S;
        S_RUN: seg_state <= SEG_C;
        S_PAUSE: seg_state <= SEG_P;
        S_ERROR: seg_state <= SEG_E;
        default: seg_state <= SEG_BLANK;
    endcase
end

// ========== ��� ==========
assign LG1 = seg_state;

// ========== �Ż�����ʾ�߼� ==========
// �ж��Ƿ���ʾ����ֵ������״̬������ɣ��������С���ͣ������״̬�µ�����ɣ�

// ��������
always @( posedge clk ) begin
     
    if( state == S_SETUP ) begin
        LG2 <= light_state ? pills_ones : 4'b0000;  // ��λ
        LG3 <= light_state ? pills_tens : 4'b0000;  // ʮλ

        LG4 <= light_state ? total_ones : 4'b0000;  // ��λ
        LG5 <= light_state ? total_tens : 4'b0000;  // ʮλ
        LG6 <= light_state ? total_hundreds : 4'b0000;  // ��λ
    end else begin
        LG2 <= (finished == 1'b1) ? pills_ones : current_pills_ones;  // ��λ
        LG3 <= (finished == 1'b1) ? pills_tens : current_pills_tens;  // ʮλ

        LG4 <= (finished == 1'b1) ? total_ones : done_ones;          // ��λ
        LG5 <= (finished == 1'b1) ? total_tens : done_tens;          // ʮλ
        LG6 <= (finished == 1'b1) ? total_hundreds : done_hundreds;  // ��λ
    end

end

// ========== ����������߼� ==========
// ������ģʽ�£�ʹ��500Hz�������������ݾ������࿪��/�ر�
// �����ʾ��ģʽ�£�����500Hz������
assign buzzer = (
    (beep_mode == BEEP_COMPLETE) ? (beep_enable && beep_tone) :  // �����ʾ����500Hz������
    (beep_mode == BEEP_ALARM || beep_mode == BEEP_ALARM_FAST) ? (beep_enable && alarm_enable && beep_tone) : // ��������500Hz������
    1'b0
);

endmodule