module clock(
    input clk,           // 1000Hz��ʱ���ź�
    input set_clr,       // ��������������ģʽ����ʱ��ͣ
    input set_clk,       // ������ѡ�е����ּ�һ
    input set_hour,      // ������ѡ������Сʱģʽ��ǰ���ǽ�������ģʽ
    input set_min,       // ������ѡ�����÷���ģʽ��ǰ���ǽ�������ģʽ
    input set_sec,       // ������ѡ��������ģʽ��ǰ���ǽ�������ģʽ
    input rst,           // ��������λ�����㿪ʼ��ʱ
    output [6:0] seg,    // ���λ���߶�����������
    output [3:0] sec,    // ��ʮλ
    output [3:0] thi,    // �ָ�λ
    output [3:0] four,   // ��ʮλ
    output [3:0] five,   // ʱ��λ
    output [3:0] six     // ʱʮλ
);

// ����������
reg [3:0] cnt;        // ���λ������
reg [3:0] sec_cnt;    // ��ʮλ������
reg [3:0] thi_cnt;    // �ָ�λ������
reg [3:0] four_cnt;   // ��ʮλ������
reg [3:0] five_cnt;   // ʱ��λ������
reg [3:0] six_cnt;    // ʱʮλ������

// ��Ƶ��������1000Hz -> 1Hz��
reg [9:0] clk_div_cnt; // 0~999������10λ�㹻����1000��
wire clk_1hz;          // 1Hz�봥���ź�

// ����������
reg set_clk_prev;     // ���ڼ��set_clk��������
wire set_clk_rise;    // set_clk�������ź�

// ---------------------- 1. 1000Hz -> 1Hz ��Ƶ�߼� ----------------------
always @(posedge clk or negedge rst) begin
    if (!rst) begin
        clk_div_cnt <= 10'b0000000000;
    end else begin
        // ������999��1000�Σ������㣬����1Hz����
        if (clk_div_cnt == 10'b1111100111) begin // 999
            clk_div_cnt <= 10'b0000000000;
        end else begin
            clk_div_cnt <= clk_div_cnt + 10'b0000000001;
        end
    end
end
// ����Ƶ��������999ʱ��clk_1hz����һ��ʱ�����ڵĸߵ�ƽ��1ms��
assign clk_1hz = (clk_div_cnt == 10'b1111100111) ? 1'b1 : 1'b0;

// ---------------------- 2. set_clk���������ؼ�⣨1000Hz������ ----------------------
always @(posedge clk or negedge rst) begin
    if (!rst) begin
        set_clk_prev <= 1'b0;
    end else begin
        set_clk_prev <= set_clk;
    end
end
assign set_clk_rise = set_clk & ~set_clk_prev;

// ---------------------- 3. ��λ�ͼ�ʱ/����ģʽ�߼� ----------------------
always @(posedge clk or negedge rst) begin
    if (!rst) begin
        // ��λ���м�����
        cnt <= 4'b0000;
        sec_cnt <= 4'b0000;
        thi_cnt <= 4'b0000;
        four_cnt <= 4'b0000;
        five_cnt <= 4'b0000;
        six_cnt <= 4'b0000;
    end else if (set_clr) begin
        // ����ģʽ����������ʱѡ��λ��1��1000Hz��ⰴ�������ӳ٣�
        if (set_clk_rise) begin
            if (set_hour) begin
                // ����Сʱ��24Сʱ�Ʊ߽紦��
                if (five_cnt == 4'b1001) begin
                    five_cnt <= 4'b0000;
                    if (six_cnt == 4'b0010) begin
                        six_cnt <= 4'b0000;
                    end else begin
                        six_cnt <= six_cnt + 4'b0001;
                    end
                end else if (six_cnt == 4'b0010 && five_cnt == 4'b0011) begin
                    // 23���ص�00��
                    five_cnt <= 4'b0000;
                    six_cnt <= 4'b0000;
                end else begin
                    five_cnt <= five_cnt + 4'b0001;
                end
            end else if (set_min) begin
                // ���÷��ӣ�60���ӱ߽紦��
                if (thi_cnt == 4'b1001) begin
                    thi_cnt <= 4'b0000;
                    if (four_cnt == 4'b0101) begin
                        four_cnt <= 4'b0000;
                    end else begin
                        four_cnt <= four_cnt + 4'b0001;
                    end
                end else begin
                    thi_cnt <= thi_cnt + 4'b0001;
                end
            end else if (set_sec) begin
                // �����루60��߽紦��
                if (cnt == 4'b1001) begin
                    cnt <= 4'b0000;
                    if (sec_cnt == 4'b0101) begin
                        sec_cnt <= 4'b0000;
                    end else begin
                        sec_cnt <= sec_cnt + 4'b0001;
                    end
                end else begin
                    cnt <= cnt + 4'b0001;
                end
            end
        end
    end else begin
        // ������ʱģʽ������1Hz�����崥��ʱ��λ
        if (clk_1hz) begin
            // ���λ������0~9��
            if (cnt == 4'b1001) begin
                cnt <= 4'b0000;
                // ��ʮλ������0~5��
                if (sec_cnt == 4'b0101) begin
                    sec_cnt <= 4'b0000;
                    // �ָ�λ������0~9��
                    if (thi_cnt == 4'b1001) begin
                        thi_cnt <= 4'b0000;
                        // ��ʮλ������0~5��
                        if (four_cnt == 4'b0101) begin
                            four_cnt <= 4'b0000;
                            // ʱ��λ+ʱʮλ������24Сʱ�ƣ�
                            if (six_cnt == 4'b0010 && five_cnt == 4'b0011) begin
                                // 23:59:59 -> 00:00:00
                                five_cnt <= 4'b0000;
                                six_cnt <= 4'b0000;
                            end else if (five_cnt == 4'b1001) begin
                                five_cnt <= 4'b0000;
                                six_cnt <= six_cnt + 4'b0001;
                            end else begin
                                five_cnt <= five_cnt + 4'b0001;
                            end
                        end else begin
                            four_cnt <= four_cnt + 4'b0001;
                        end
                    end else begin
                        thi_cnt <= thi_cnt + 4'b0001;
                    end
                end else begin
                    sec_cnt <= sec_cnt + 4'b0001;
                end
            end else begin
                cnt <= cnt + 4'b0001;
            end
        end
    end
end

// ---------------------- 4. �߶������������ ----------------------
reg [6:0] seg_out;
always @(*) begin
    case(cnt)
        4'b0000: seg_out = 7'b0111111;  // ��ʾ����0
        4'b0001: seg_out = 7'b0000110;  // ��ʾ����1
        4'b0010: seg_out = 7'b1011011;  // ��ʾ����2
        4'b0011: seg_out = 7'b1001111;  // ��ʾ����3
        4'b0100: seg_out = 7'b1100110;  // ��ʾ����4
        4'b0101: seg_out = 7'b1101101;  // ��ʾ����5
        4'b0110: seg_out = 7'b1111101;  // ��ʾ����6
        4'b0111: seg_out = 7'b0000111;  // ��ʾ����7
        4'b1000: seg_out = 7'b1111111;  // ��ʾ����8
        4'b1001: seg_out = 7'b1101111;  // ��ʾ����9
        default: seg_out = 7'b0000000; // Ĭ��Ϩ��
    endcase
end

// �����ֵ
assign seg = seg_out;
assign sec = sec_cnt;
assign thi = thi_cnt;
assign four = four_cnt;
assign five = five_cnt;
assign six = six_cnt;

endmodule