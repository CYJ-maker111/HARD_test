module clock(
    input clk,           // 1000Hz��ʱ���ź�
    input set_clr,       // ��������������ģʽ����ʱ��ͣ
    input set_clk,       // ������ѡ�е����ּ�һ
    input set_hour,      // ������ѡ������Сʱģʽ��ǰ���ǽ�������ģʽ
    input set_min,       // ������ѡ�����÷���ģʽ��ǰ���ǽ�������ģʽ
    input set_sec,       // ������ѡ��������ģʽ��ǰ���ǽ�������ģʽ
    input rst,           // ��������λ�����㿪ʼ��ʱ
    output [6:0] seg,    // ���λ���߶�����������
    output [3:0] sec,    // ��ʮλ
    output [3:0] thi,    // �ָ�λ
    output [3:0] four,   // ��ʮλ
    output [3:0] five,   // ʱ��λ
    output [3:0] six     // ʱʮλ
);

// ����������
reg [3:0] cnt;        // ���λ������
reg [3:0] sec_cnt;    // ��ʮλ������
reg [3:0] thi_cnt;    // �ָ�λ������
reg [3:0] four_cnt;   // ��ʮλ������
reg [3:0] five_cnt;   // ʱ��λ������
reg [3:0] six_cnt;    // ʱʮλ������

// ��Ƶ��������1000Hz -> 1Hz��
reg [9:0] clk_div_cnt; // 0~999������10λ�㹻����1000��
wire clk_1hz;          // 1Hz�봥���ź�

// ����������
reg set_clk_prev;     // ���ڼ��set_clk��������
wire set_clk_rise;    // set_clk�������ź�

// ʱ�䳣�����壨�����ɶ��ԣ�
localparam MAX_SEC_ONES  = 4'b1001; // ���λ���ֵ9
localparam MAX_SEC_TENS  = 4'b0101; // ��ʮλ���ֵ5
localparam MAX_MIN_ONES  = 4'b1001; // �ָ�λ���ֵ9
localparam MAX_MIN_TENS  = 4'b0101; // ��ʮλ���ֵ5
localparam MAX_HOUR_ONES = 4'b1001; // ʱ��λ���ֵ9
localparam MAX_HOUR_TENS = 4'b0010; // ʱʮλ���ֵ2
localparam HOUR_23_ONES  = 4'b0011; // 23ʱ�ĸ�λ3

// ����������������ģʽ��ѡ���ź�תΪ��ֵ������case��
reg [1:0] set_mode;
always @(*) begin
    if (set_sec)      set_mode = 2'b01; // ������
    else if (set_min) set_mode = 2'b10; // ���÷�
    else if (set_hour)set_mode = 2'b11; // ����ʱ
    else              set_mode = 2'b00; // ��ѡ��
end

// ---------------------- 1. 1000Hz -> 1Hz ��Ƶ�߼� ----------------------
always @(posedge clk or negedge rst) begin
    if (!rst) begin
        clk_div_cnt <= 10'b0000000000;
    end else begin
        if (clk_div_cnt == 10'b1111100111) begin // 999
            clk_div_cnt <= 10'b0000000000;
        end else begin
            clk_div_cnt <= clk_div_cnt + 10'b0000000001;
        end
    end
end
assign clk_1hz = (clk_div_cnt == 10'b1111100111) ? 1'b1 : 1'b0;

// ---------------------- 2. set_clk���������ؼ�� ----------------------
always @(posedge clk or negedge rst) begin
    if (!rst) begin
        set_clk_prev <= 1'b0;
    end else begin
        set_clk_prev <= set_clk;
    end
end
assign set_clk_rise = set_clk & ~set_clk_prev;

// ---------------------- 3. ����ʱ/�����߼����޸�23:59:59��λ�� ----------------------
always @(posedge clk or negedge rst) begin
    if (!rst) begin
        // ��λ���м�����
        cnt <= 4'b0000;
        sec_cnt <= 4'b0000;
        thi_cnt <= 4'b0000;
        four_cnt <= 4'b0000;
        five_cnt <= 4'b0000;
        six_cnt <= 4'b0000;
    end 
    // ģʽ1������ģʽ����������ʱ�䣬��case���if-else if��
    else if (set_clr && set_clk_rise) begin
        case(set_mode)
            2'b01: begin // ������
                if (cnt == MAX_SEC_ONES) begin
                    cnt <= 4'b0000;
                    sec_cnt <= (sec_cnt == MAX_SEC_TENS) ? 4'b0000 : (sec_cnt + 4'b0001);
                end else begin
                    cnt <= cnt + 4'b0001;
                end
            end
            2'b10: begin // ���÷�
                if (thi_cnt == MAX_MIN_ONES) begin
                    thi_cnt <= 4'b0000;
                    four_cnt <= (four_cnt == MAX_MIN_TENS) ? 4'b0000 : (four_cnt + 4'b0001);
                end else begin
                    thi_cnt <= thi_cnt + 4'b0001;
                end
            end
            2'b11: begin // ����ʱ
                if (six_cnt == MAX_HOUR_TENS && five_cnt == HOUR_23_ONES) begin
                    five_cnt <= 4'b0000;
                    six_cnt <= 4'b0000;
                end else if (five_cnt == MAX_HOUR_ONES) begin
                    five_cnt <= 4'b0000;
                    six_cnt <= six_cnt + 4'b0001;
                end else begin
                    five_cnt <= five_cnt + 4'b0001;
                end
            end
            default: ; // ��ѡ�񣬲�����
        endcase
    end
    // ģʽ2��������ʱģʽ���ؼ��޸�������ʱ�߼��ж�˳��
    else if (!set_clr && clk_1hz) begin
        // ---------------------- �롢�ֽ�λ�߼���ԭ�߼����䣩 ----------------------
        // ����1�����λ��λ��9��0��
        if (cnt == MAX_SEC_ONES) begin
            cnt <= 4'b0000;
        end else begin
            cnt <= cnt + 4'b0001;
        end
        // ����2����ʮλ��λ��59���0�룩
        if (cnt == MAX_SEC_ONES && sec_cnt == MAX_SEC_TENS) begin
            sec_cnt <= 4'b0000;
        end else if (cnt == MAX_SEC_ONES) begin
            sec_cnt <= sec_cnt + 4'b0001;
        end
        // ����3���ָ�λ��λ��59�����+1��9��0��
        if (cnt == MAX_SEC_ONES && sec_cnt == MAX_SEC_TENS && thi_cnt == MAX_MIN_ONES) begin
            thi_cnt <= 4'b0000;
        end else if (cnt == MAX_SEC_ONES && sec_cnt == MAX_SEC_TENS) begin
            thi_cnt <= thi_cnt + 4'b0001;
        end
        // ����4����ʮλ��λ��59�֡�0�֣�
        if (cnt == MAX_SEC_ONES && sec_cnt == MAX_SEC_TENS && thi_cnt == MAX_MIN_ONES && four_cnt == MAX_MIN_TENS) begin
            four_cnt <= 4'b0000;
        end else if (cnt == MAX_SEC_ONES && sec_cnt == MAX_SEC_TENS && thi_cnt == MAX_MIN_ONES) begin
            four_cnt <= four_cnt + 4'b0001;
        end

        // ---------------------- ʱ��λ�߼��������޸��������ж�˳�� ----------------------
        // �����ȼ���ߡ�����5��23:59:59 �� 00:00:00 ȫ������
        if (cnt == MAX_SEC_ONES && sec_cnt == MAX_SEC_TENS && thi_cnt == MAX_MIN_ONES && four_cnt == MAX_MIN_TENS 
            && six_cnt == MAX_HOUR_TENS && five_cnt == HOUR_23_ONES) begin
            five_cnt <= 4'b0000;
            six_cnt <= 4'b0000;
        end
        // ����6��ʱ��λ��9��ʱʮλ��1���� 09:59:59 �� 10:00:00��
        else if (cnt == MAX_SEC_ONES && sec_cnt == MAX_SEC_TENS && thi_cnt == MAX_MIN_ONES && four_cnt == MAX_MIN_TENS 
                && five_cnt == MAX_HOUR_ONES) begin
            five_cnt <= 4'b0000;
            six_cnt <= six_cnt + 4'b0001;
        end
        // ����7����ͨ�����ʱ��λ��1���� 12:59:59 �� 13:00:00��
        else if (cnt == MAX_SEC_ONES && sec_cnt == MAX_SEC_TENS && thi_cnt == MAX_MIN_ONES && four_cnt == MAX_MIN_TENS) begin
            five_cnt <= five_cnt + 4'b0001;
        end
    end
end

// ---------------------- 4. �߶������������ ----------------------
reg [6:0] seg_out;
always @(*) begin
    case(cnt)
        4'b0000: seg_out = 7'b0111111;  // ��ʾ����0
        4'b0001: seg_out = 7'b0000110;  // ��ʾ����1
        4'b0010: seg_out = 7'b1011011;  // ��ʾ����2
        4'b0011: seg_out = 7'b1001111;  // ��ʾ����3
        4'b0100: seg_out = 7'b1100110;  // ��ʾ����4
        4'b0101: seg_out = 7'b1101101;  // ��ʾ����5
        4'b0110: seg_out = 7'b1111101;  // ��ʾ����6
        4'b0111: seg_out = 7'b0000111;  // ��ʾ����7
        4'b1000: seg_out = 7'b1111111;  // ��ʾ����8
        4'b1001: seg_out = 7'b1101111;  // ��ʾ����9
        default: seg_out = 7'b0000000; // Ĭ��Ϩ��
    endcase
end

// �����ֵ
assign seg = seg_out;
assign sec = sec_cnt;
assign thi = thi_cnt;
assign four = four_cnt;
assign five = five_cnt;
assign six = six_cnt;

endmodule